-- format_leaf.vhd
-- $ : Log
-- @ : Author
-- # : Section
-- % : Outer interface
-- ! : Caution!
-- ? : Question
-- & :
-- * :
-- + :
-- ^ :
-- | :
-- () :
-- [] :
-- {} :

